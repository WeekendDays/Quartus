LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY led2 IS
PORT(a7: IN STD_LOGIC;
	 x7: OUT STD_LOGIC);
END led2;

ARCHITECTURE led2a OF led2 IS
BEGIN
	x7 <= a7;
END led2a;