LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mydecoder3_8_1 IS
	PORT(a: in STD_LOGIC_VECTOR(2 DOWNTO 0);
		 d: out STD_LOGIC_VECTOR(7 DOWNTO 0));
END mydecoder3_8_1;

ARCHITECTURE decoder OF mydecoder3_8_1 IS
BEGIN
	d <= "10000000" WHEN a = "000" ELSE
		 "01000000" WHEN a = "001" ELSE
		 "00100000" WHEN a = "010" ELSE
		 "00010000" WHEN a = "011" ELSE
		 "00001000" WHEN a = "100" ELSE
		 "00000100" WHEN a = "101" ELSE
		 "00000010" WHEN a = "110" ELSE
		 "00000001";
END decoder;